-----------------------------------------------------------------------
-- Multiplication and division with subroutines (divmul.asm)
-----------------------------------------------------------------------
LIBRARY ieee, work; USE ieee.std_logic_1164.ALL, work.support.ALL;
PACKAGE firmware IS
CONSTANT DefaultFrequency : DECIHERTZ := 15; -- 1 to 1000
CONSTANT SimDIP : WORD := "00000000"; -- DIP input for testbench only
CONSTANT Firmware : WORDx256  := (
0   => "00001110", 1   => "00101000",  -- CALL 40
2   => "11100000",                     -- PUSH R0
3   => "00001110", 4   => "00000111",  -- CALL 7
5   => "11110010",                     -- POP R2
6   => "00000000",                     -- HLT
7   => "00010000", 8   => "00000000",  -- MOV R0, 0
9   => "00010011", 10  => "00000001",  -- MOV R3, 1
11  => "00010001", 12  => "10110011",  -- MOV R1, 179
13  => "00010010", 14  => "00001100",  -- MOV R2, 12
15  => "00001010", 16  => "00011001",  -- JS 25
17  => "10111000", 18  => "00100001",  -- CMP R2, R1
19  => "00000100", 20  => "00011001",  -- JC 25
21  => "10100011",                     -- LSHIFT R3
22  => "10100010",                     -- LSHIFT R2
23  => "00000010", 24  => "00001111",  -- JMP 15
25  => "10111000", 26  => "00010010",  -- CMP R1, R2
27  => "00000101", 28  => "00100001",  -- JNC 33
29  => "00111000", 30  => "00010010",  -- SUB R1, R2
31  => "01011000", 32  => "00000011",  -- OR R0, R3
33  => "11010010",                     -- RSHIFT R2
34  => "11010011",                     -- RSHIFT R3
35  => "00000110", 36  => "00100111",  -- JZ 39
37  => "00000010", 38  => "00011001",  -- JMP 25
39  => "00001111",                     -- RETURN
40  => "00010000", 41  => "00000000",  -- MOV R0, 0
42  => "10010001", 43  => "01100100",  -- LOAD R1, [100]
44  => "10010010", 45  => "01100101",  -- LOAD R2, [101]
46  => "00000110", 47  => "00111010",  -- JZ 58
48  => "11000010", 49  => "00000001",  -- BIT R2, 1
50  => "00000110", 51  => "00110110",  -- JZ 54
52  => "00101000", 53  => "00000001",  -- ADD R0, R1
54  => "10100001",                     -- LSHIFT R1
55  => "11010010",                     -- RSHIFT R2
56  => "00000010", 57  => "00101110",  -- JMP 46
58  => "00001111",                     -- RETURN
100 => "00000111",                     -- 7
101 => "00011101",                     -- 29
OTHERS => "UUUUUUUU");END;