-----------------------------------------------------------------------
-- LED Matrix display test -- fills matrices 3 and 4 with counters
-----------------------------------------------------------------------
LIBRARY ieee, work; USE ieee.std_logic_1164.ALL, work.support.ALL;
PACKAGE firmware IS
CONSTANT SimDIP : WORD := "00000000";
CONSTANT InitSpeed : NATURAL := 5;
CONSTANT Firmware : WORDx256  := (
0   => "00010000", 1   => "11001000",  -- 10C8  MOV R0, 200 (-56)
2   => "00010001", 3   => "00000000",  -- 1100  MOV R1, 0
4   => "10110000", 5   => "11111111",  -- B0FF  CMP R0, 255 (-1)
6   => "00000110", 7   => "00011110",  -- 061E  JZ 30
8   => "10001000", 9   => "00010000",  -- 8810  STORE R1, [R0]
10  => "10110000", 11  => "11001111",  -- B0CF  CMP R0, 207 (-49)
12  => "00000110", 13  => "00011010",  -- 061A  JZ 26
14  => "00100000", 15  => "00000001",  -- 2001  ADD R0, 1
16  => "00000010", 17  => "00000100",  -- 0204  JMP 4
18  => "10110000", 19  => "11010000",  -- B0D0  CMP R0, 208 (-48)
20  => "00000110", 21  => "00011010",  -- 061A  JZ 26
22  => "00100000", 23  => "00000001",  -- 2001  ADD R0, 1
24  => "00000010", 25  => "00000100",  -- 0204  JMP 4
26  => "00010000", 27  => "11111000",  -- 10F8  MOV R0, 248 (-8)
28  => "00000010", 29  => "00000100",  -- 0204  JMP 4
30  => "00100001", 31  => "00000001",  -- 2101  ADD R1, 1
32  => "00010000", 33  => "11001000",  -- 10C8  MOV R0, 200 (-56)
34  => "00000010", 35  => "00000100",  -- 0204  JMP 4
OTHERS => "UUUUUUUU");END;