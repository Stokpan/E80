-----------------------------------------------------------------------
-- Olimex GateMateA1-EVB Board Settings for the E80 Computer
-- Copyright (C) 2026 Panos Stokas <panos.stokas@hotmail.com>
-----------------------------------------------------------------------
PACKAGE Board IS
CONSTANT BoardCLK_MHz : NATURAL := 10;
END;