-----------------------------------------------------------------------
-- Multiplication and division with subroutines (divmul.asm)
-----------------------------------------------------------------------
LIBRARY ieee, work; USE ieee.std_logic_1164.ALL, work.support.ALL;
PACKAGE firmware IS
CONSTANT DefaultFrequency : DECIHERTZ := 15; -- 1 to 1000
CONSTANT SimDIP : WORD := "00000000"; -- DIP input for testbench only
CONSTANT Firmware : WORDx256  := (
0   => "00001110", 1   => "00101010",  -- CALL 42
2   => "11100000",                     -- PUSH R0
3   => "00001110", 4   => "00000111",  -- CALL 7
5   => "11110010",                     -- POP R2
6   => "00000000",                     -- HLT
7   => "00010001", 8   => "10110011",  -- MOV R1, 179
9   => "00010010", 10  => "00001100",  -- MOV R2, 12
11  => "00010000", 12  => "00000000",  -- MOV R0, 0
13  => "00010011", 14  => "00000001",  -- MOV R3, 1
15  => "10111000", 16  => "00100001",  -- CMP R2, R1
17  => "00000100", 18  => "00011011",  -- JC 27
19  => "11010010", 20  => "10000000",  -- BIT R2, 128
21  => "00000111", 22  => "00011011",  -- JNZ 27
23  => "11000010",                     -- LSHIFT R2
24  => "11000011",                     -- LSHIFT R3
25  => "00000010", 26  => "00001111",  -- JMP 15
27  => "10111000", 28  => "00010010",  -- CMP R1, R2
29  => "00000101", 30  => "00100011",  -- JNC 35
31  => "00111000", 32  => "00010010",  -- SUB R1, R2
33  => "01101000", 34  => "00000011",  -- OR R0, R3
35  => "10100010",                     -- RSHIFT R2
36  => "10100011",                     -- RSHIFT R3
37  => "00000110", 38  => "00101001",  -- JZ 41
39  => "00000010", 40  => "00011011",  -- JMP 27
41  => "00001111",                     -- RETURN
42  => "10010001", 43  => "01100100",  -- LOAD R1, [100]
44  => "10010010", 45  => "01100101",  -- LOAD R2, [101]
46  => "00010000", 47  => "00000000",  -- MOV R0, 0
48  => "11010010", 49  => "11111111",  -- BIT R2, 255
50  => "00000110", 51  => "00111110",  -- JZ 62
52  => "11010010", 53  => "00000001",  -- BIT R2, 1
54  => "00000110", 55  => "00111010",  -- JZ 58
56  => "00101000", 57  => "00000001",  -- ADD R0, R1
58  => "11000001",                     -- LSHIFT R1
59  => "10100010",                     -- RSHIFT R2
60  => "00000010", 61  => "00110000",  -- JMP 48
62  => "00001111",                     -- RETURN
100 => "00000111",                     -- 7
101 => "00011101",                     -- 29
OTHERS => "UUUUUUUU");END;