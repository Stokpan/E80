-----------------------------------------------------------------------
-- DivMul.e80asm - Unsigned division and multiplication
-----------------------------------------------------------------------
LIBRARY ieee, work; USE ieee.std_logic_1164.ALL, work.support.ALL;
PACKAGE firmware IS
CONSTANT SimDIP : WORD := "00000000";
CONSTANT InitSpeed : NATURAL := 4;
CONSTANT Firmware : WORDx256  := (
0   => "00001110", 1   => "00101000",  -- 0E28  CALL 40
2   => "11100000",                     -- E0    PUSH R0
3   => "00001110", 4   => "00000111",  -- 0E07  CALL 7
5   => "11110010",                     -- F2    POP R2
6   => "00000000",                     -- 00    HLT
7   => "00010000", 8   => "00000000",  -- 1000  MOV R0, 0
9   => "00010011", 10  => "00000001",  -- 1301  MOV R3, 1
11  => "00010001", 12  => "10110011",  -- 11B3  MOV R1, 179 (-77)
13  => "00010010", 14  => "00001100",  -- 120C  MOV R2, 12
15  => "00001010", 16  => "00011001",  -- 0A19  JS 25
17  => "10111000", 18  => "00100001",  -- B821  CMP R2, R1
19  => "00000100", 20  => "00011001",  -- 0419  JC 25
21  => "10100011",                     -- A3    LSHIFT R3
22  => "10100010",                     -- A2    LSHIFT R2
23  => "00000010", 24  => "00001111",  -- 020F  JMP 15
25  => "10111000", 26  => "00010010",  -- B812  CMP R1, R2
27  => "00000101", 28  => "00100001",  -- 0521  JNC 33
29  => "00111000", 30  => "00010010",  -- 3812  SUB R1, R2
31  => "01011000", 32  => "00000011",  -- 5803  OR R0, R3
33  => "11010010",                     -- D2    RSHIFT R2
34  => "11010011",                     -- D3    RSHIFT R3
35  => "00000110", 36  => "00100111",  -- 0627  JZ 39
37  => "00000010", 38  => "00011001",  -- 0219  JMP 25
39  => "00001111",                     -- 0F    RETURN
40  => "00010000", 41  => "00000000",  -- 1000  MOV R0, 0
42  => "00010001", 43  => "00000111",  -- 1107  MOV R1, 7
44  => "00010010", 45  => "00011101",  -- 121D  MOV R2, 29
46  => "00000110", 47  => "00111010",  -- 063A  JZ 58
48  => "11000010", 49  => "00000001",  -- C201  BIT R2, 1
50  => "00000110", 51  => "00110110",  -- 0636  JZ 54
52  => "00101000", 53  => "00000001",  -- 2801  ADD R0, R1
54  => "10100001",                     -- A1    LSHIFT R1
55  => "11010010",                     -- D2    RSHIFT R2
56  => "00000010", 57  => "00101110",  -- 022E  JMP 46
58  => "00001111",                     -- 0F    RETURN
OTHERS => "UUUUUUUU");END;